module singleseconds (reset, clk, enable, ss, nxt);
  input reset, clk, enable;
  output [3:0] ss;
  output       nxt;
  reg    [3:0] ss;
  
  assign nxt= (ss == 4'd9);
  always @(posedge clk or posedge reset)
    if (reset) ss <= 4'd0;
      else if (enable)
             if (nxt) ss <= 0;
               else ss <= ss + 1;
endmodule



module tenthsofseconds (reset, clk, enable, ts);
  input reset, clk, enable;
  output [2:0] ts;
  wire         again;
  reg    [2:0] ts;
  
  assign again = (ts == 3'd5);
  always @(posedge clk or posedge reset)
    if (reset) ts <= 4'd0;
      else if (enable)
             if (again) ts <= 0;
               else ts <= ts + 1;
endmodule



module secondcounter (reset, clk, enable, enablet, ts, ss, st);
  input reset, clk, enable, enablet;
  output [2:0] ts;
  output [3:0] ss;
  output [3:0] st;
  wire         ent, ens;

  
  singleseconds   i0 (reset, clk, enable & ens, ss, ent);
  tenthsofseconds i1 (reset, clk, enable & ent, ts);
  singleseconds	atenth	(reset, clk, enablet, st, ens);

endmodule


/*
module test();
  reg reset, clk;
  wire [2:0] ts;
  wire [3:0] ss;

  secondcounter CUT (reset, clk, 1'b1, ts, ss);
  
  initial begin reset =0; clk = 0; #10 reset = 1; #9 reset = 0; end
  always #4 clk = ~clk;
endmodule
*/