`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:  University of Patras
// Engineer: iTalos
// 
// Create Date:    15:41:27 09/25/2023 
// Design Name: 
// Module Name:    Character_Memory 
// Project Name:   iTalos
//
//////////////////////////////////////////////////////////////////////////////////
module Character_Memory(
	 input Pixelclock,
    input [7:0] character,
    output [8:0] RGB
    );
	 
	 reg memory_counter [
	 


endmodule
